
--
--  Consolidated Data Load script for odbcapture_installation_logs data
--
--  Must be run as SYSTEM
--
--  Command Line Parameters:
--   1 - SYSTEM/password@TNSALIAS
--       i.e. pass the username and password for the SYSTEM user
--            and the TNSALIAS for the connection to the database.
--       The Data Load installation requires this connection information.
--

prompt
prompt Confirm/Create odbcapture_installation_logs Table
declare
   jnk  number := 0;
   procedure run_sql (in_sql in varchar2) is begin
      dbms_output.put_line(in_sql || ';');
      execute immediate in_sql;
   exception when others then
      dbms_output.put_line('-- ' || SQLERRM || CHR(10));
   end run_sql;
begin
   begin
      execute immediate 'insert into odbcapture_installation_logs(load_dtm, install_type, file_name)' ||
                        ' values(sysdate, ''Test'', ''Test'')';
      rollback;
      jnk := 1;
   exception when others then
      if SQLERRM != 'ORA-00942: table or view does not exist'
      then
         dbms_output.put_line('odbcapture_installation_logs table: ' || SQLERRM);
      end if;
      jnk := -1;
   end;
   if jnk = -1
   then
      run_sql('create table odbcapture_installation_logs' || CHR(10) ||
         ' (load_dtm date' || CHR(10) ||
         ' ,install_type varchar2(10)' || CHR(10) ||
         ' ,file_name varchar2(512)' || CHR(10) ||
         ' ,contents clob)');
      run_sql('comment on column odbcapture_installation_logs.load_dtm is ''Date/Time the installation log file was loaded.''');
      run_sql('comment on column odbcapture_installation_logs.install_type is ''Type of installation (from TYPE_CONF).''');
      run_sql('comment on column odbcapture_installation_logs.file_name is ''Name of installation log file.''');
      run_sql('comment on column odbcapture_installation_logs.contents is ''Contents/Text of the installation log file.''');
      run_sql('comment on table odbcapture_installation_logs is ''ODBCAPTURE installation log files.''');
      run_sql('grant select on odbcapture_installation_logs to public');
      run_sql('create public synonym odbcapture_installation_logs for odbcapture_installation_logs');
   end if;
end;
/


-- NOTE: Additional file extensions for SQL*Loader include
--   .bad - Bad Records
--   .dsc - Discard Records
--   .log - Log File

prompt
prompt sqlldr_control=./odbcapture_installation_logs.ctl
host sqlldr '&1.' control=odbcapture_installation_logs.ctl data=odbcapture_installation_logs.csv log=odbcapture_installation_logs.log silent=HEADER,FEEDBACK

begin
   if '&_RC.' != '0' then
      raise_application_error(-20000, 'Control file "odbcapture_installation_logs.ctl" returned error: &_RC.');
   end if;
end;
/

